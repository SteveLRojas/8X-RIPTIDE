library verilog;
use verilog.vl_types.all;
entity hazard_unit is
    port(
        clk             : in     vl_logic;
        NZT1            : in     vl_logic;
        NZT2            : in     vl_logic;
        NZT3            : in     vl_logic;
        NZT4            : in     vl_logic;
        JMP             : in     vl_logic;
        XEC1            : in     vl_logic;
        XEC2            : in     vl_logic;
        XEC3            : in     vl_logic;
        XEC4            : in     vl_logic;
        RET             : in     vl_logic;
        CALL4           : in     vl_logic;
        ALU_NZ          : in     vl_logic;
        alu_op          : in     vl_logic_vector(2 downto 0);
        alu_mux         : in     vl_logic;
        HALT            : in     vl_logic;
        RST             : in     vl_logic;
        regf_a_read     : in     vl_logic_vector(2 downto 0);
        regf_w_reg1     : in     vl_logic_vector(2 downto 0);
        regf_w_reg2     : in     vl_logic_vector(2 downto 0);
        regf_w_reg3     : in     vl_logic_vector(2 downto 0);
        regf_w_reg4     : in     vl_logic_vector(2 downto 0);
        regf_w_reg5     : in     vl_logic_vector(2 downto 0);
        regf_wren_reg1  : in     vl_logic;
        regf_wren_reg2  : in     vl_logic;
        regf_wren_reg3  : in     vl_logic;
        regf_wren_reg4  : in     vl_logic;
        regf_wren_reg5  : in     vl_logic;
        SC_reg1         : in     vl_logic;
        SC_reg2         : in     vl_logic;
        SC_reg3         : in     vl_logic;
        SC_reg4         : in     vl_logic;
        SC_reg5         : in     vl_logic;
        SC_reg6         : in     vl_logic;
        SC_reg7         : in     vl_logic;
        WC_reg1         : in     vl_logic;
        WC_reg2         : in     vl_logic;
        WC_reg3         : in     vl_logic;
        WC_reg4         : in     vl_logic;
        WC_reg5         : in     vl_logic;
        WC_reg6         : in     vl_logic;
        WC_reg7         : in     vl_logic;
        n_LB_w_reg1     : in     vl_logic;
        n_LB_w_reg2     : in     vl_logic;
        n_LB_w_reg3     : in     vl_logic;
        n_LB_w_reg4     : in     vl_logic;
        n_LB_w_reg5     : in     vl_logic;
        n_LB_w_reg6     : in     vl_logic;
        n_LB_w_reg7     : in     vl_logic;
        n_LB_r          : in     vl_logic;
        rotate_mux      : in     vl_logic;
        rotate_source   : in     vl_logic;
        latch_wren      : in     vl_logic;
        latch_wren1     : in     vl_logic;
        latch_wren2     : in     vl_logic;
        latch_address_w1: in     vl_logic_vector(1 downto 0);
        latch_address_w2: in     vl_logic_vector(1 downto 0);
        latch_address_r : in     vl_logic_vector(1 downto 0);
        shift_L         : in     vl_logic_vector(2 downto 0);
        hazard          : out    vl_logic;
        branch_hazard   : out    vl_logic;
        pipeline_flush  : out    vl_logic;
        decoder_RST     : out    vl_logic
    );
end hazard_unit;
